`timescale 1ns / 1ps

module RST_SYNC_tb ();

/////////////////////////////////////////////////////
//////////////////clk_generator//////////////////////
/////////////////////////////////////////////////////

parameter clk_period= 20; 
reg clk_tb=0; 
always #(clk_period/2) clk_tb = ~clk_tb;

/////////////////////////////////////////////////////
///////////////Decleration & Instances///////////////
/////////////////////////////////////////////////////

reg       rst_tb;
wire      sync_rst_tb;

 RST_SYNC DUT (
		.clk(clk_tb),
		.rst(rst_tb),
		.sync_rst(sync_rst_tb)
		);


/////////////////////////////////////////////////////
///////////////////Initial Block/////////////////////
/////////////////////////////////////////////////////

initial begin 
	$dumpfile("BIT_SYNC.vcd"); 
	$dumpvars; 
	
	reset();
	
end 

/////////////////////////////////////////////////////
//////////////////////Tasks//////////////////////////
/////////////////////////////////////////////////////

task reset;
 begin
 rst_tb=1;
 #(clk_period)
 rst_tb=0;
 #(clk_period)
 rst_tb=1;
 end
endtask

endmodule
