`timescale 1ns / 1ps

module BIT_SYNC_tb ();

parameter BUS_WIDTH = 5 ;

/////////////////////////////////////////////////////
//////////////////clk_generator//////////////////////
/////////////////////////////////////////////////////
parameter clk_period= 20; 
reg clk_tb=0; 
always #(clk_period/2) clk_tb = ~clk_tb;

/////////////////////////////////////////////////////
///////////////Decleration & Instances///////////////
/////////////////////////////////////////////////////

reg	[BUS_WIDTH - 1:0]       	async_tb;
reg		                        rst_tb;
wire [BUS_WIDTH - 1:0]			sync_tb;

 BIT_SYNC #(BUS_WIDTH) DUT (
		.async(async_tb),
		.clk(clk_tb),
		.rst(rst_tb),
		.sync(sync_tb)
		);


/////////////////////////////////////////////////////
///////////////////Initial Block/////////////////////
/////////////////////////////////////////////////////

initial begin 
	$dumpfile("BIT_SYNC.vcd"); 
	$dumpvars; 
	
	reset();
	
	async_tb = 5'b10101;
end 

/////////////////////////////////////////////////////
//////////////////////Tasks//////////////////////////
/////////////////////////////////////////////////////

task reset;
 begin
 rst_tb=1;
 #(clk_period)
 rst_tb=0;
 #(clk_period)
 rst_tb=1;
 end
endtask
endmodule
